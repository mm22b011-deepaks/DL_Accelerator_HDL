`define STATE_DIM 4
`define MAT_DIM 4

