`define MAT_DIM 4
`define bits_int 16
`define bits_frac 16
